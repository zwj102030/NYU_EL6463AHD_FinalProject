----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    15:34:27 11/13/2017
-- Design Name:
-- Module Name:    DataMemory - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
--Library work;
use work.def.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DataMemory is
    Port ( Address : in  STD_LOGIC_VECTOR (31 downto 0);
           WrtData : in  STD_LOGIC_VECTOR (31 downto 0);
           clk : in  STD_LOGIC;
           we : in  STD_LOGIC;
			  ukey : in  STD_LOGIC_VECTOR (127 downto 0);
			  Din : in  STD_LOGIC_VECTOR (63 downto 0);
           RdData : out  STD_LOGIC_VECTOR (31 downto 0);
			  Dout : out  STD_LOGIC_VECTOR (63 downto 0);
			  en_din : in  STD_LOGIC;
			  en_ukey : in  STD_LOGIC;
			  clr : in  STD_LOGIC;
			  RAM_OUT : out RAM_Array);
end DataMemory;

architecture Behavioral of DataMemory is

--type RAM_Array is array (0 to 63) --This is 10000 x 32bits RAM
--	of std_logic_vector(31 downto 0);
signal RAM : RAM_array:=
( 0 => "10110111111000010101000101100011",
1 => "01010110000110001100101100011100",
2 => "11110100010100000100010011010101",
3 => "10010010100001111011111010001110",
4 => "00110000101111110011100001000111",
5 => "11001110111101101011001000000000",
6 => "01101101001011100010101110111001",
7 => "00001011011001011010010101110010",
8 => "10101001100111010001111100101011",
9 => "01000111110101001001100011100100",
10 => "11100110000011000001001010011101",
11 => "10000100010000111000110001010110",
12 => "00100010011110110000011000001111",
13 => "11000000101100100111111111001000",
14 => "01011110111010011111100110000001",
15 => "11111101001000010111001100111010",
16 => "10011011010110001110110011110011",
17 => "00111001100100000110011010101100",
18 => "11010111110001111110000001100101",
19 => "01110101111111110101101000011110",
20 => "00010100001101101101001111010111",
21 => "10110010011011100100110110010000",
22 => "01010000101001011100011101001001",
23 => "11101110110111010100000100000010",
24 => "10001101000101001011101010111011",
25 => "00101011010011000011010001110100",
26 => x"a1b2a1b2",
27 => x"3333a1b2", 
28 => x"3333a1b2", 
29 => x"a1b2a1b2", 
30 => x"a1b2abab",
31 => x"a1b2ee88",

 others => (others=>'0') );

begin
	
	Process1 :process(clk)
		begin
		
		if( en_din = '1' or en_ukey = '1')then
					RAM(26) <= ukey( 127 downto 96);
					RAM(27) <= ukey( 95 downto 64);
					RAM(28) <= ukey( 63 downto 32);
					RAM(29) <= ukey( 31 downto 0);
					RAM(30) <= Din( 63 downto 32);
					RAM(31) <= Din( 31 downto 0);
		end if;
		
      -- RESET
			if (clr = '1') then
				RAM(0) <= "10110111111000010101000101100011";
				RAM(1) <= "01010110000110001100101100011100";
				RAM(2) <= "11110100010100000100010011010101";
				RAM(3) <= "10010010100001111011111010001110";
				RAM(4) <= "00110000101111110011100001000111";
				RAM(5) <= "11001110111101101011001000000000";
				RAM(6) <= "01101101001011100010101110111001";
				RAM(7) <= "00001011011001011010010101110010";
				RAM(8) <= "10101001100111010001111100101011";
				RAM(9) <= "01000111110101001001100011100100";
				RAM(10) <= "11100110000011000001001010011101";
				RAM(11) <= "10000100010000111000110001010110";
				RAM(12) <= "00100010011110110000011000001111";
				RAM(13) <= "11000000101100100111111111001000";
				RAM(14) <= "01011110111010011111100110000001";
				RAM(15) <= "11111101001000010111001100111010";
				RAM(16) <= "10011011010110001110110011110011";
				RAM(17) <= "00111001100100000110011010101100";
				RAM(18) <= "11010111110001111110000001100101";
				RAM(19) <= "01110101111111110101101000011110";
				RAM(20) <= "00010100001101101101001111010111";
				RAM(21) <= "10110010011011100100110110010000";
				RAM(22) <= "01010000101001011100011101001001";
				RAM(23) <= "11101110110111010100000100000010";
				RAM(24) <= "10001101000101001011101010111011";
				RAM(25) <= "00101011010011000011010001110100";
				------
					RAM(26) <= ukey( 127 downto 96);
					RAM(27) <= ukey( 95 downto 64);
					RAM(28) <= ukey( 63 downto 32);
					RAM(29) <= ukey( 31 downto 0);
					RAM(30) <= Din( 63 downto 32);
					RAM(31) <= Din( 31 downto 0);
--				RAM(26) <= x"00000000";
--				RAM(27) <= x"00000000";
--				RAM(28) <= x"00000000";
--				RAM(29) <= x"00000000";
--				RAM(30) <= x"00000000";
--				RAM(31) <= x"00000000";
--				RAM(32) <= x"00000000";
--				RAM(33) <= x"00000000";
--				RAM(34) <= x"00000000";
--				RAM(35) <= x"00000000";
--				RAM(36) <= x"00000000";
--				RAM(37) <= x"00000000";
--				RAM(38) <= x"00000000";
--				RAM(39) <= x"00000000";
--				RAM(40) <= x"00000000";
--				RAM(41) <= x"00000000";
--				RAM(42) <= x"00000000";
--				RAM(43) <= x"00000000";
--				RAM(44) <= x"00000000";
--				RAM(45) <= x"00000000";
--				RAM(46) <= x"00000000";
--				RAM(47) <= x"00000000";
--				RAM(48) <= x"00000000";
--				RAM(49) <= x"00000000";
--				RAM(50) <= x"00000000";
--				RAM(51) <= x"00000000";
--				RAM(52) <= x"00000000";
--				RAM(53) <= x"00000000";
--				RAM(54) <= x"00000000";
--				RAM(55) <= x"00000000";
--				RAM(56) <= x"00000000";
--				RAM(57) <= x"00000000";
--				RAM(58) <= x"00000000";
--				RAM(59) <= x"00000000";
--				RAM(60) <= x"00000000";
--				RAM(61) <= x"00000000";
--				RAM(62) <= x"00000000";
--				RAM(63) <= x"00000000";
					--RAM(31) <= Din( 31 downto 0);
			elsif (clk = '1' and clk'Event) then
				if we = '1' then


					RAM(conv_integer('0'&Address(5 downto 0))) <= WrtData;
				--else RdData <= RAM(conv_integer(Address));
				end if;

--				if en_ukey = '1' then
-----------------------------------------------------------------------------------------------------------------------
--          RAM(0) <= "10110111111000010101000101100011";
--          RAM(1) <= "01010110000110001100101100011100";
--          RAM(2) <= "11110100010100000100010011010101";
--          RAM(3) <= "10010010100001111011111010001110";
--          RAM(4) <= "00110000101111110011100001000111";
--          RAM(5) <= "11001110111101101011001000000000";
--          RAM(6) <= "01101101001011100010101110111001";
--          RAM(7) <= "00001011011001011010010101110010";
--          RAM(8) <= "10101001100111010001111100101011";
--          RAM(9) <= "01000111110101001001100011100100";
--          RAM(10) <= "11100110000011000001001010011101";
--          RAM(11) <= "10000100010000111000110001010110";
--          RAM(12) <= "00100010011110110000011000001111";
--          RAM(13) <= "11000000101100100111111111001000";
--          RAM(14) <= "01011110111010011111100110000001";
--          RAM(15) <= "11111101001000010111001100111010";
--          RAM(16) <= "10011011010110001110110011110011";
--          RAM(17) <= "00111001100100000110011010101100";
--          RAM(18) <= "11010111110001111110000001100101";
--          RAM(19) <= "01110101111111110101101000011110";
--          RAM(20) <= "00010100001101101101001111010111";
--          RAM(21) <= "10110010011011100100110110010000";
--          RAM(22) <= "01010000101001011100011101001001";
--          RAM(23) <= "11101110110111010100000100000010";
--          RAM(24) <= "10001101000101001011101010111011";
--          RAM(25) <= "00101011010011000011010001110100";
-----------------------------------------------------------------------------------------------------------------------
--					RAM(26) <= ukey( 127 downto 96);
--					RAM(27) <= ukey( 95 downto 64);
--					RAM(28) <= ukey( 63 downto 32);
--					RAM(29) <= ukey( 31 downto 0);
--				end if;
--
--				if en_din = '1' then
--					RAM(30) <= x"FFFFFFFF";---Din( 63 downto 32);
--					RAM(31) <= Din( 31 downto 0);
--				end if;
			end if;
		end process;

	with we select RdData <=
	    RAM(conv_integer('0'&Address(5 downto 0))) when '0',
		 x"00000000" when others;

	Dout <= RAM(32) & RAM(33);
	RAM_OUT <= RAM;

end Behavioral;
