----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    19:14:22 11/10/2017
-- Design Name:
-- Module Name:    ROM_2to32_32bit - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM_2to32_32bit is
    Port ( Address : in  STD_LOGIC_VECTOR (31 downto 0);
           Data : out  STD_LOGIC_VECTOR (31 downto 0));
end ROM_2to32_32bit;

architecture Behavioral of ROM_2to32_32bit is

type ROM_Array is array (0 to 400) --This is 10000 x 32bits ROM

	of std_logic_vector(31 downto 0);

--Suppose ROM has been prestored value like this table
    constant Content: ROM_Array := (

--	 --test 1:
--        0 => "00000000000000000000000000000000",		-- in dian's design, this instruction is ignored;
--        1 => "00001100000000010000000000000000",		-- ANDI: R1 = R0 &(000...0), i.e. R1=0;
--        2 => "00000000001000010000000000010000",		-- ADD: R0=R1+R1, i.e. R0=0;
--        3 => "00000100000000010001000100100010",      -- ADDI: R1=R0+signext(1122)=1122(hex), R0=0;
--        4 => "00000100000000000001000100010001",		-- ADDI: R0=R0+1111=1111(hex);
--        5 => "00000000001000000001000000010001",      -- SUB: R2=R1-R0=0011(hex), R1=1122,R0=1111,R2=0011;
--        6 => "00001000000000110000000000010001",      -- SUBI: R3=R0-0011=1100(hex), R0 checked;
--		  7 => "00000000001000110010000000010010",      -- AND: R4=R1&R3=1122&1100=1100(hex);
--		  8 => "00000000001000100010100000010011",      -- OR: R5=R1|R2=1122|0011=1133(hex), R1,R2 checked;
--		  9 => "00010000001001100100011100000000",      -- ORI: R6=R1|4700=1122|4700=5722(hex), R1 checked;
--		  10 => "00000000001000110011100000010100",     -- NOR: R7=!(R1|R3)=11111111111111111110111011011101, R3 checked;
--		  11 => "00000000100001010100000000010000",     -- ADD: R8=R4+R5,check R4, R5;
--		 -- 12 => "11111100110001110000000000000000",     -- HALT: STOP & check R6, R7;
--
--
--	 --test 2: SW & LW
--	     12 => "00100000010000010000000000000001",     -- SW: R1 -> MEM[0011+1],i.e. MEM[0012]=1122;
--	     13 => "00100000000001100001000100010001",     -- SW: R6 -> MEM[1111+1111], i.e. MEM[2222]=5722;
--		  14 => "00011100010000110000000000000001",     -- LW: MEM[0011+1] -> R3, i.e. R3=1122;
--        15 => "00011101010001000010001000100010",     -- LW: MEM[0+2222] -> R4, i.e. R4=5722;
--		  16 => "00000000100000111000000000010000",		-- ADD: R16=R4+R3, i.e. Rs:R4,Rt:R3, check R4,R3; (checked)
--	--	  17 => "11111100000000000000000000000000",     -- HALT: STOP ;
--
--
--	--test 4: SHL & SHR
--		  17 => "00010100011010000000000000000100",		-- SHL: R8=R3<<<imm(4), i.e. R8=R3<<<4; R8=11220
--		  18 => "00011000100001110000000000000011",		-- SHR: R7=R4>>>imm(3), i.e. R7=R4>>>3; R7=ae4
--		  19 => "11111100111010000000000000000000",     -- HALT: STOP ; check R7,R8 (checked)
--
--		  20 => "00000100000000010001000100100010",
--		  21 => "00000000100000111000000000010000",
--		  22 => "11111100111010000000000000000000",


-- --key_exp
"00000000000000000000000000000000", -- 0
"00000100000000010000000000000000", ---1
"00000100000000100000000000000000",---2
"00000100000000110000000000000000",---3
"00000100000001000000000000000000",---4
"00000100000001010000000000000000",----5
"00000100000001100000000000000000",----6
"00000100000001110000000000000000",---7
"00000100000010000000000000000000",---8
"00000100000010010000000000000000",----9
"00000100000010100000000000000000",---10
"00000100000010110000000000000000",---11
"00000100000011000000000000000000",---12
"00000100000011010000000000000000",----13
"00000100000011100000000000000000",---14
"00000100000011110000000000000000",----15
"00000100000100000000000000000000",----16
"00000100000100010000000000000000",-----17
"00000100000100100000000000000000",----18
"00000100000100110000000000000000",---19
"00000100000000010000000000000000", -- 1 start of key_exp
"00101100000000001111111111111111", -- BNE R0 R0 -1
"00000100000000100000000000000000",
"00000100000000110000000000000000",
"00000100000010000000000000000100",
"00000100000010010000000001001110",
"00000100000001000000000000011010",
"00101100100000100000000000000001",
"00000100000000100000000000000000",
"00101101000000110000000000000001",
"00000100000000110000000000000000",
"00011100010001100000000000000000",
"00000001010010110110000000010000",
"00000001100001100110100000010000",
"00010101101011000000000000000011",
"00011001101011100000000000011101",
"00000001100011100110100000010011",
"00100000010011010000000000000000",
"00000101101010100000000000000000",
"00011100011001010000000000011010",
"00000001010010110110000000010000",
"00000001100001010110100000010000",
"00101001100000000000000000000110",
"00010101101011100000000000000001",
"00011001101011110000000000011111",
"00000001110011110110100000010011",
"00001001100011110000000000000001",
"00001101111011000000000000011111",
"00101101100000001111111111111010",
"00100000011011010000000000011010",
"00000101101010110000000000000000",
"00000100010001110000000000000001",
"00000100111000100000000000000000",
"00000100011001110000000000000001",
"00000100111000110000000000000000",
"00000100001001110000000000000001",
"00000100111000010000000000000000",
"00101100001010011111111111100000",
"00101000000000001111111111111111", --38 end of key_exp
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000", --100
"00001100000000000000000000000000", -- 101 start of enc
"00001100001000010000000000000000",
"00001100010000100000000000000000",
"00001100011000110000000000000000",
"00001100100001000000000000000000",
"00001100101001010000000000000000",
"00001100110001100000000000000000",
"00001100111001110000000000000000",
"00001101000010000000000000000000",
"00001101001010010000000000000000",
"00001101010010100000000000000000",
"00001101011010110000000000000000",
"00001101100011000000000000000000",
"00001101101011010000000000000000",
"00001101110011100000000000000000",
"00001101111011110000000000000000",
"00001110000100000000000000000000",
"00001110001100010000000000000000",
"00001110010100100000000000000000",
"00001110011100110000000000000000",
"00001110100101000000000000000000",
"00011100000000100000000000011110",
"00011100000000110000000000011111",
"00000100101001010000000000001101",
"00000100110001100000000000000001",
"00000110011100110000000000000001",
"00010110011100110000000000011111",
"00000110010100100000000000011111",
"00011100000000010000000000000000",
"00000000001000100001000000010000",
"00011100110001110000000000000000",
"00000000111000110001100000010000",
"00000010010000111010000000010010",
"00000000010000110100100000010010",
"00000000010000110101000000010100",
"00000001001010100100000000010100",
"00101010100000000000000000000110",
"00000010011010000101100000010010",
"00010101000010000000000000000001",
"00000101100011000000000000000001",
"00101001011000000000000000000001",
"00000101000010000000000000000001",
"00101101100101001111111111111010",
"00010100110011100000000000000001",
"00011101110011110000000000000000",
"00000001111010000001000000010000",
"00000010010000101010000000010010",
"00000000010000110100100000010010",
"00000000010000110101000000010100",
"00000001001010100100000000010100",
"00000100000011000000000000000000",
"00101010100000000000000000000110",
"00000010011010000101100000010010",
"00010101000010000000000000000001",
"00000101100011000000000000000001",
"00101001011000000000000000000001",
"00000101000010000000000000000001",
"00101101100101001111111111111010",
"00000101110100000000000000000001",
"00011101110100010000000000000001",
"00000010001010000001100000010000",
"00000100110001100000000000000001",
"00000100000011000000000000000000",
"00101100110001011111111111100000",
"00100000000000100000000000100000",
"00100000000000110000000000100001",
"00101000000000001111111111111111", --end of enc
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000", --200
"00001100000000000000000000000000",
"00001100001000010000000000000000",
"00001100010000100000000000000000",
"00001100011000110000000000000000",
"00001100100001000000000000000000",
"00001100101001010000000000000000",
"00001100110001100000000000000000",
"00001100111001110000000000000000",
"00001101000010000000000000000000",
"00001101001010010000000000000000",
"00001101010010100000000000000000",
"00001101011010110000000000000000",
"00001101100011000000000000000000",
"00001101101011010000000000000000",
"00001101110011100000000000000000",
"00001101111011110000000000000000",
"00001110000100000000000000000000",
"00001110001100010000000000000000",
"00001110010100100000000000000000",
"00001110011100110000000000000000",
"00001110100101000000000000000000",
"00011100000001010000000000011110",
"00011100000001100000000000011111",
"00000100001000010000000000001100",
"00000100000000100000000000000001",
"00010100010100110000000000011111",
"00000110010100100000000000011111",
"00010100001000110000000000000001",
"00000010010001011010000000010010",
"00011100011001000000000000000001",
"00000000110001000011100000010001",
"00101010100000000000000000000110",
"00000000010001110100000000010010",
"00011000111001110000000000000001",
"00000101001010010000000000000001",
"00101001000000000000000000000001",
"00000000111100110011100000010000",
"00101101001101001111111111111001",
"00000000111001010101000000010010",
"00000000111001010101100000010100",
"00000001010010110011000000010100",
"00000010010001101010000000010010",
"00000100000010010000000000000000",
"00011100011011000000000000000000",
"00000000101011000011100000010001",
"00101010100000000000000000000110",
"00000000010001110100000000010010",
"00011000111001110000000000000001",
"00000101001010010000000000000001",
"00101001000000000000000000000001",
"00000000111100110011100000010000",
"00101101001101001111111111111001",
"00000100000010010000000000000000",
"00000000111001100101000000010010",
"00000000111001100101100000010100",
"00000001010010110010100000010100",
"00001000001000010000000000000001",
"00101100001000001111111111100001",
"00000101101011010000000000000001",
"00011100000011100000000000000001",
"00011100000011110000000000000000",
"00000000110011101000000000010001",
"00000000101011111000100000010001",
"00100000000100010000000000100010",
"00100000000100000000000000100011",
"00101000000000001111111111111111", --end of dec


		OTHERS => "00000000000000000000000000000000"
	);
begin
	process1: process(Address)
	begin
		Data <= Content(conv_integer(Address(9 downto 0)));
	end process;

end Behavioral;
